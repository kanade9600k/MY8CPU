/* Tennis game Program */
// テニスゲームのプログラム
module ROM_B(address, data);

input [7:0] address;
output [15:0] data;

wire [7:0] address;
reg [15:0] data;

always @* begin
    
    case (address)
        8'b00000000: data <= 16'b00100010_10000000; // MOV A, 128
        8'b00000001: data <= 16'b00101100_00000000; // OUT A
        8'b00000010: data <= 16'b00000010_00000000; // ADD A, 0 タイミング調整
        8'b00000011: data <= 16'b00101001_00000000; // IN B
        8'b00000100: data <= 16'b00001011_00000011; // AND B, 3
        8'b00000101: data <= 16'b00000011_11111101; // ADD B, 253
        8'b00000110: data <= 16'b00110000_00110111; // JNC 55 ノーマルモードのスタートにジャンプ
        8'b00000111: data <= 16'b00011100_00000000; // SR A ハードモードスタート地点
        8'b00001000: data <= 16'b00111100_11111010; // SET C, 250
        8'b00001001: data <= 16'b00101100_00000000; // OUT A
        8'b00001010: data <= 16'b00000010_00000000; // ADD A, 0 タイミング調整
        8'b00001011: data <= 16'b00000010_00000000; // ADD A, 0 タイミング調整
        8'b00001100: data <= 16'b00101001_00000000; // IN B 一番外の無限ループスタート地点 □ ■
        8'b00001101: data <= 16'b00001011_00000001; // AND B, 1
        8'b00001110: data <= 16'b00000011_11111111; // ADD B, 255
        8'b00001111: data <= 16'b00110000_00010101; // JNC 21 終了処理の下のアドレスまでジャンプ
        8'b00010000: data <= 16'b00100010_00000000; // MOV A, 0 左勝利の終了処理開始
        8'b00010001: data <= 16'b00101100_00000000; // OUT A
        8'b00010010: data <= 16'b00100010_11110000; // MOV A, 240
        8'b00010011: data <= 16'b00101100_00000000; // OUT A
        8'b00010100: data <= 16'b00110100_00110110; // JMP 54 プログラム終了のアドレスまでジャンプ
        8'b00010101: data <= 16'b00011100_00000000; // SR A スルーしたときはここにジャンプ
        8'b00010110: data <= 16'b00101100_00000000; // OUT A
        8'b00010111: data <= 16'b00111000_00000001; // INC C, 1
        8'b00011000: data <= 16'b00110000_00001100; // JNC 12 ループ終了点 ■
        8'b00011001: data <= 16'b00101001_00000000; // IN B 
        8'b00011010: data <= 16'b00001011_00000001; // AND B, 1
        8'b00011011: data <= 16'b00000011_11111111; // ADD B, 255
        8'b00011100: data <= 16'b00110000_00010000; // JNC 16 0なら左勝利の終了処理開始までジャンプ
        8'b00011101: data <= 16'b00011000_00000000; // SL A
        8'b00011110: data <= 16'b00101100_00000000; // OUT A
        8'b00011111: data <= 16'b00111100_11111010; // SET C, 250
        8'b00100000: data <= 16'b00000010_00000000; // ADD A, 0 タイミング調整
        8'b00100001: data <= 16'b00101001_00000000; // IN B ループ開始点 ■
        8'b00100010: data <= 16'b00001011_00000010; // AND B, 2
        8'b00100011: data <= 16'b00000011_11111111; // ADD B, 255
        8'b00100100: data <= 16'b00110000_00101010; // JNC 42 終了処理の下のアドレスまでジャンプ
        8'b00100101: data <= 16'b00100010_00000000; // MOV A, 0  右勝利の終了処理開始
        8'b00100110: data <= 16'b00101100_00000000; // OUT A
        8'b00100111: data <= 16'b00100010_00001111; // MOV A, 15
        8'b00101000: data <= 16'b00101100_00000000; // OUT A
        8'b00101001: data <= 16'b00110100_00110110; // JMP 54 プログラム終了のアドレス 
        8'b00101010: data <= 16'b00011000_00000000; // SL A スルーしたときはここにジャンプ
        8'b00101011: data <= 16'b00101100_00000000; // OUT A
        8'b00101100: data <= 16'b00111000_00000001; // INC C, 1
        8'b00101101: data <= 16'b00110000_00100001; // JNC 33 ループ終了点 ■
        8'b00101110: data <= 16'b00101001_00000000; // IN B 
        8'b00101111: data <= 16'b00001011_00000010; // AND B, 2
        8'b00110000: data <= 16'b00000011_11111111; // ADD B, 255
        8'b00110001: data <= 16'b00110000_00100101; // JNC 37 0なら右勝利の終了処理開始までジャンプ
        8'b00110010: data <= 16'b00011100_00000000; // SR A
        8'b00110011: data <= 16'b00101100_00000000; // OUT A
        8'b00110100: data <= 16'b00111100_11111010; // SET C, 250
        8'b00110101: data <= 16'b00110100_00001100; // JMP 12 無限ループの終了点 □
        8'b00110110: data <= 16'b00110100_00110110; // JMP 54 自分自身にジャンプ(プログラム終了) *****プログラムの終了地点*****
        // この下から編集
        8'b00110111: data <= 16'b00000010_00000000; // ノーマルモードスタート地点 タイミング調整
        8'b00111000: data <= 16'b00000010_00000000; // ADD A, 0タイミング調整
        8'b00111001: data <= 16'b00000010_00000000; // ADD A, 0タイミング調整
        8'b00111010: data <= 16'b00000010_00000000; // ADD A, 0タイミング調整
        8'b00111011: data <= 16'b00000010_00000000; // ADD A, 0タイミング調整
        8'b00111100: data <= 16'b00011100_00000000; // SR A 
        8'b00111101: data <= 16'b00111100_11111010; // SET C, 250
        8'b00111110: data <= 16'b00101100_00000000; // OUT A
        8'b00111111: data <= 16'b00000010_00000000; // ADD A, 0 タイミング調整
        8'b01000000: data <= 16'b00000010_00000000; // ADD A, 0 タイミング調整
        8'b01000001: data <= 16'b00101001_00000000; // IN B 一番外の無限ループスタート地点 □ ■
        8'b01000010: data <= 16'b00001011_00000001; // AND B, 1
        8'b01000011: data <= 16'b00000011_11111111; // ADD B, 255
        8'b01000100: data <= 16'b00110000_01001010; // JNC 74 終了処理の下のアドレスまでジャンプ
        8'b01000101: data <= 16'b00100010_00000000; // MOV A, 0 左勝利の終了処理開始
        8'b01000110: data <= 16'b00101100_00000000; // OUT A
        8'b01000111: data <= 16'b00100010_11110000; // MOV A, 240
        8'b01001000: data <= 16'b00101100_00000000; // OUT A
        8'b01001001: data <= 16'b00110100_00110110; // JMP 54 プログラム終了のアドレスまでジャンプ
        8'b01001010: data <= 16'b00011100_00000000; // SR A スルーしたときはここにジャンプ
        8'b01001011: data <= 16'b00000010_00000000; // ADD A, 0タイミング調整
        8'b01001100: data <= 16'b00000010_00000000; // ADD A, 0タイミング調整
        8'b01001101: data <= 16'b00000010_00000000; // ADD A, 0タイミング調整
        8'b01001110: data <= 16'b00000010_00000000; // ADD A, 0タイミング調整
        8'b01001111: data <= 16'b00000010_00000000; // ADD A, 0タイミング調整
        8'b01010000: data <= 16'b00101100_00000000; // OUT A
        8'b01010001: data <= 16'b00111000_00000001; // INC C, 1
        8'b01010010: data <= 16'b00110000_01000001; // JNC 65 ループ終了点 ■
        8'b01010011: data <= 16'b00000010_00000000; // ADD A, 0タイミング調整
        8'b01010100: data <= 16'b00000010_00000000; // ADD A, 0タイミング調整
        8'b01010101: data <= 16'b00000010_00000000; // ADD A, 0タイミング調整
        8'b01010110: data <= 16'b00000010_00000000; // ADD A, 0タイミング調整
        8'b01010111: data <= 16'b00000010_00000000; // ADD A, 0タイミング調整
        8'b01011000: data <= 16'b00101001_00000000; // IN B 
        8'b01011001: data <= 16'b00001011_00000001; // AND B, 1
        8'b01011010: data <= 16'b00000011_11111111; // ADD B, 255
        8'b01011011: data <= 16'b00110000_01000101; // JNC 69 0なら左勝利の終了処理開始までジャンプ
        8'b01011100: data <= 16'b00011000_00000000; // SL A
        8'b01011101: data <= 16'b00101100_00000000; // OUT A
        8'b01011110: data <= 16'b00111100_11111010; // SET C, 250
        8'b01011111: data <= 16'b00000010_00000000; // ADD A, 0 タイミング調整
        8'b01100000: data <= 16'b00101001_00000000; // IN B ループ開始点 ■
        8'b01100001: data <= 16'b00001011_00000010; // AND B, 2
        8'b01100010: data <= 16'b00000011_11111111; // ADD B, 255
        8'b01100011: data <= 16'b00110000_01101001; // JNC 105 終了処理の下のアドレスまでジャンプ
        8'b01100100: data <= 16'b00100010_00000000; // MOV A, 0  右勝利の終了処理開始
        8'b01100101: data <= 16'b00101100_00000000; // OUT A
        8'b01100110: data <= 16'b00100010_00001111; // MOV A, 15
        8'b01100111: data <= 16'b00101100_00000000; // OUT A
        8'b01101000: data <= 16'b00110100_00110110; // JMP 54 プログラム終了のアドレス 
        8'b01101001: data <= 16'b00011000_00000000; // SL A スルーしたときはここにジャンプ
        8'b01101010: data <= 16'b00000010_00000000; // ADD A, 0タイミング調整
        8'b01101011: data <= 16'b00000010_00000000; // ADD A, 0タイミング調整
        8'b01101100: data <= 16'b00000010_00000000; // ADD A, 0タイミング調整
        8'b01101101: data <= 16'b00000010_00000000; // ADD A, 0タイミング調整
        8'b01101110: data <= 16'b00000010_00000000; // ADD A, 0タイミング調整
        8'b01101111: data <= 16'b00101100_00000000; // OUT A
        8'b01110000: data <= 16'b00111000_00000001; // INC C, 1
        8'b01110001: data <= 16'b00110000_01100000; // JNC 96 ループ終了点 ■
        8'b01110010: data <= 16'b00000010_00000000; // ADD A, 0タイミング調整
        8'b01110011: data <= 16'b00000010_00000000; // ADD A, 0タイミング調整
        8'b01110100: data <= 16'b00000010_00000000; // ADD A, 0タイミング調整
        8'b01110101: data <= 16'b00000010_00000000; // ADD A, 0タイミング調整
        8'b01110110: data <= 16'b00000010_00000000; // ADD A, 0タイミング調整
        8'b01110111: data <= 16'b00101001_00000000; // IN B 
        8'b01111000: data <= 16'b00001011_00000010; // AND B, 2
        8'b01111001: data <= 16'b00000011_11111111; // ADD B, 255
        8'b01111010: data <= 16'b00110000_01100100; // JNC 100 0なら右勝利の終了処理開始までジャンプ
        8'b01111011: data <= 16'b00011100_00000000; // SR A
        8'b01111100: data <= 16'b00101100_00000000; // OUT A
        8'b01111101: data <= 16'b00111100_11111010; // SET C, 250
        8'b01111110: data <= 16'b00110100_01000001; // JMP 65 無限ループの終了点 □
        default: data <= 16'bxxxxxxxx_xxxxxxxx;
    endcase
end

endmodule